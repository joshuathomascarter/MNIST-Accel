/*
  systolic_array.v - Weight-Stationary Systolic Array
  ---------------------------------------------------
  ARCHITECTURAL CORRECTION:
   - This is a WEIGHT-STATIONARY (WS) array.
   - Weights are broadcast to columns and stored in PEs.
   - Activations stream horizontally (West -> East).
   - Partial sums accumulate locally in each PE.
   
  Engineer's Note:
   - This module instantiates an NxM grid of PEs.
   - The 'row_en' signal is critical for power gating unused rows during
     sparse operations or small matrix multiplications.
   - Ensure 'load_weight' is asserted for at least 1 cycle before 'en' goes high.
   
  Parameters:
   N_ROWS : number of rows (default 2)
   N_COLS : number of columns (default 2)
   PIPE   : pass to each PE (1 inserts internal pipeline)
   SAT    : pass to each mac8 instance inside PE
   ENABLE_CLOCK_GATING: 1 enables BUFGCE/ICG insertion for power savings.
*/
`ifndef SYSTOLIC_ARRAY_V
`define SYSTOLIC_ARRAY_V
`default_nettype none
// -----------------------------------------------------------------------------
// Title      : systolic_array
// File       : systolic_array.v
// Description: Weight-Stationary INT8 systolic array with Pk=1.
//              Verilog-2001 compliant; uses generate loops and flattened ports.
//
//              WEIGHT-STATIONARY DATAFLOW:
//              - Weights loaded ONCE and stored stationary in each PE
//              - Activations stream horizontally (west to east)
//              - No vertical weight flow (weights broadcast to all PEs in same column)
//              - Maximum weight reuse efficiency
//
// Requirements Trace:
//   REQ-ACCEL-SYST-01: Provide N_ROWS x N_COLS grid of PEs accumulating INT32 psums.
//   REQ-ACCEL-SYST-02: Stream activations (A) from west edge, broadcast weights (B) to columns.
//   REQ-ACCEL-SYST-03: Support synchronous clear of all partial sums via clr.
//   REQ-ACCEL-SYST-04: Deterministic hold when en=0.
//   REQ-ACCEL-SYST-05: Support weight preloading via load_weight control.
//   REQ-ACCEL-SYST-06: Optional single-cycle pipeline inside each PE (PIPE param).
// -----------------------------------------------------------------------------
// Parameters:
//   N_ROWS : number of rows (default 2)
//   N_COLS : number of columns (default 2)
//   PIPE   : pass to each PE (1 inserts internal pipeline)
//   SAT    : pass to each mac8 instance inside PE
// -----------------------------------------------------------------------------
// Port Flattening:
//   a_in_flat  [N_ROWS*8-1:0] contains N_ROWS signed 8-bit lanes (row-major)
//   b_in_flat  [N_COLS*8-1:0] contains N_COLS signed 8-bit lanes (col-major)
//   c_out_flat [N_ROWS*N_COLS*32-1:0] concatenated row-major
//   load_weight: when high, PEs capture b_in and store stationary
// -----------------------------------------------------------------------------
module systolic_array #(
  parameter N_ROWS = 14,
  parameter N_COLS = 14,
  parameter PIPE   = 1,
  parameter ENABLE_CLOCK_GATING = 1
)(
  input  wire clk,
  input  wire rst_n,
  input  wire en,
  input  wire clr,
  input  wire load_weight,
  input  wire [N_ROWS-1:0] row_en,
  input  wire [N_ROWS*N_COLS-1:0] bypass_flat,  // ← ADD THIS: Per-PE bypass signal
  input  wire [N_ROWS*8-1:0] a_in_flat,
  input  wire [N_COLS*8-1:0] b_in_flat,
  output wire [N_ROWS*N_COLS*32-1:0] c_out_flat
);

  // ---------------------------------------------------------------------------
  // 1. Input Unpacking & SKEW GENERATION (Triangular Shift Register)
  // ---------------------------------------------------------------------------
  
  wire signed [7:0] a_in_raw [0:N_ROWS-1]; // Raw inputs from flat bus
  wire signed [7:0] a_in     [0:N_ROWS-1]; // Skewed inputs to array
  wire signed [7:0] b_in     [0:N_COLS-1];

  genvar ui;
  generate
    // Unpack raw inputs
    for (ui = 0; ui < N_ROWS; ui = ui + 1) begin : UNPACK_A_RAW
      assign a_in_raw[ui] = a_in_flat[ui*8 +: 8];
    end
    
    // Unpack weights (No skew needed for broadcast weights in WS)
    for (ui = 0; ui < N_COLS; ui = ui + 1) begin : UNPACK_B
      assign b_in[ui] = b_in_flat[ui*8 +: 8];
    end
    
    // NEW: Unpack bypass signals (Per-PE bypass for residual connections in ResNet)
    for (ui = 0; ui < N_ROWS*N_COLS; ui = ui + 1) begin : UNPACK_BYPASS
      integer r_idx, c_idx;
      initial begin
        r_idx = ui / N_COLS;
        c_idx = ui % N_COLS;
      end
      assign bypass_mat[r_idx][c_idx] = bypass_flat[ui];
    end

    // Create Triangular Skew for Activations
    // Row 0: 0 delays
    // Row 1: 1 delay
    // ...
    // Row N: N delays
    for (ui = 0; ui < N_ROWS; ui = ui + 1) 
    
      if (ui == 0) begin
        // Row 0 goes straight through
        assign a_in[ui] = a_in_raw[ui];
      end else begin
        // Rows 1..N get shift registers
        reg signed [7:0] delay_regs [0:ui-1]; // Array of registers of size 'ui'
        integer k;
        
        always @(posedge clk or negedge rst_n) begin
          if (!rst_n) begin
            for (k=0; k<ui; k=k+1) delay_regs[k] <= 8'sd0;
          end else if (en) begin
            // Shift register logic
            delay_regs[0] <= a_in_raw[ui];
            for (k=1; k<ui; k=k+1) begin
               delay_regs[k] <= delay_regs[k-1];
            end
          end
        end
        assign a_in[ui] = delay_regs[ui-1]; // Output of the last delay register
      end
  
  endgenerate

  // ========================================================================
  // 2. Clock Gating (Per-Row) - Saves 434 mW @ 100 MHz
  // ========================================================================
  // Engineer's Note:
  // This is a critical power optimization. By gating the clock to unused rows,
  // we eliminate dynamic power consumption in the PEs (which are the main consumers).
  // When ENABLE_CLOCK_GATING=1, each row gets gated clock (gates when !row_en[i])
  // When ENABLE_CLOCK_GATING=0, all rows use main clock (for simulation/debug)
  // Uses Xilinx BUFGCE primitive for glitch-free clock gating
  
  wire [N_ROWS-1:0] row_clk;  // Gated clocks per row
  
  generate
    if (ENABLE_CLOCK_GATING) begin : gen_clock_gating
      for (ui = 0; ui < N_ROWS; ui = ui + 1) begin : gen_row_gates
        wire row_clk_en;
        // CRITICAL FIX: Clock must be active for Compute (en), Weight Load (load_weight), or Clear (clr)
        // Previously: assign row_clk_en = en & row_en[ui]; (This prevented weight loading!)
        assign row_clk_en = row_en[ui] & (en | load_weight | clr);
        
        // Xilinx BUFGCE: Clock buffer with gate enable (glitch-free)
        // For ASIC: use integrated clock gate cell (ICG) from library
        `ifdef XILINX_FPGA
          BUFGCE row_clk_gate (
            .I  (clk),
            .CE (row_clk_en),
            .O  (row_clk[ui])
          );
        `else
          // Generic clock gating (use latch-based gate for glitch-free operation)
          reg row_clk_en_latched;
          always @(clk or row_clk_en) begin
            if (!clk) row_clk_en_latched <= row_clk_en;  // Latch on falling edge
          end
          assign row_clk[ui] = clk & row_clk_en_latched;
        `endif
      end
    end else begin : gen_no_clock_gating
      // No clock gating - all rows use main clock
      for (ui = 0; ui < N_ROWS; ui = ui + 1) begin : gen_row_direct_clk
        assign row_clk[ui] = clk;
      end
    end
  endgenerate

  // ---------------------------------------------------------------------------
  // 3. PE Grid Instantiation
  // ---------------------------------------------------------------------------
  // Engineer's Note:
  // This double loop generates the physical grid of PEs.
  // - Activations (a_src) are chained horizontally.
  // - Weights (b_src) are BROADCAST vertically (all PEs in col 'c' get b_in[c]).
  // - This confirms the Weight-Stationary architecture.
  
  // Forwarding nets between PEs (ONLY for activations, NOT weights!)
  wire signed [7:0] a_fwd [0:N_ROWS-1][0:N_COLS-1];
  wire signed [31:0] acc_mat [0:N_ROWS-1][0:N_COLS-1];
  
  // NEW: Forwarding nets for load_weight (Systolic Fanout Fix)
  wire load_weight_fwd [0:N_ROWS-1][0:N_COLS-1];
  
  // NEW: 2D bypass matrix for residual mode (ResNet support)
  wire bypass_mat [0:N_ROWS-1][0:N_COLS-1];

  genvar r, c;
  generate
    for (r = 0; r < N_ROWS; r = r + 1) begin : ROW
      for (c = 0; c < N_COLS; c = c + 1) begin : COL
        // Activation source: from west edge or left neighbor
        wire signed [7:0] a_src = (c == 0) ? a_in[r] : a_fwd[r][c-1];
        
        // Weight source: BROADCAST from top edge to ALL rows in this column
        // NO vertical weight flow - same weight to all PEs in a column!
        wire signed [7:0] b_src = b_in[c];  // Direct from input, no forwarding
        
        // NEW: Load Weight source: From scheduler (col 0) or left neighbor
        wire load_weight_src = (c == 0) ? load_weight : load_weight_fwd[r][c-1];
        
        pe #(.PIPE(PIPE)) u_pe (
          .clk(row_clk[r]),  // Use gated clock per row
          .rst_n(rst_n),
          .a_in(a_src), 
          .b_in(b_src),  // Weight broadcast (not forwarded from neighbor)
          .bypass(bypass_mat[r][c]),  // NEW: Bypass signal for residual mode
          .en(en), 
          .clr(clr),
          .load_weight(load_weight_src),  // NEW: Chained load_weight
          .a_out(a_fwd[r][c]),
          .load_weight_out(load_weight_fwd[r][c]), // NEW: Pass to neighbor
          // b_out removed - no weight forwarding!
          .acc(acc_mat[r][c])
        );
      end
    end
  endgenerate

  // ---------------------------------------------------------------------------
  // 4. Output Packing
  // ---------------------------------------------------------------------------
  // Engineer's Note:
  // Flattens the 2D array of results into a single wide bus.
  // Uses SystemVerilog streaming operator for cleaner syntax.
  
  assign c_out_flat = { >> {acc_mat} };

  // ---------------------------------------------------------------------------
  // 5. Assertions & Verification
  // ---------------------------------------------------------------------------
  // Engineer's Note: These assertions verify the control protocol.
  
  `ifdef ASSERT_ON
    // 1. Mutual Exclusion: Cannot Compute and Load Weights simultaneously
    //    (This would corrupt the stationary weights or produce garbage psums)
    property p_mutex_load_compute;
      @(posedge clk) disable iff (!rst_n) (load_weight |-> !en);
    endproperty
    assert property (p_mutex_load_compute) 
      else $error("SYSTOLIC_ERROR: 'en' and 'load_weight' asserted simultaneously!");

    // 2. Clock Gating Safety: If we are active, ensure row_en is not all zeros
    //    (If global controls are high but all rows are disabled, we are stalling)
    property p_valid_activity;
      @(posedge clk) disable iff (!rst_n) ((en | load_weight | clr) |-> |row_en);
    endproperty
    cover property (p_valid_activity);

    // 3. Reset Check: When reset is asserted, output should eventually be 0
    //    (Note: This is a liveness property, simplified here)
    property p_reset_clears;
      @(posedge clk) !rst_n |=> (c_out_flat == 0);
    endproperty
    cover property (p_reset_clears);
  `endif

endmodule
`endif
`default_nettype wire
