/*
  mac8.v - Signed 8x8 -> 16 multiply-accumulate with 32-bit accumulator
  --------------------------------------------------------------------
  Purpose
    Small, unit-exact MAC used by the Accel v1 systolic array.  Multiplies
    two signed 8-bit inputs and accumulates into a signed 32-bit register.
    Optional saturation mode and a per-cycle saturation flag are provided.

  Key properties
    - Input:  signed [7:0] a, b
    - Product: signed [15:0] prod16 = a * b
    - Accumulator: signed [31:0] acc_r
    - Controls:
        en  : enable accumulation this cycle (when 1, compute acc := acc + a*b)
        clr : synchronous clear (when 1, acc := 0 on next clock)
        rst_n: active-low reset, clears accumulator
    - SAT parameter:
        SAT = 1 -> clamp accumulator to INT32_MIN/INT32_MAX on overflow
        SAT = 0 -> wrap-around semantics, but sat_flag still reports overflow
    - sat_flag pulses when a signed overflow/underflow is detected on the addition.

  Overflow detection (signed two's complement)
    - Signed overflow for sum = X + Y happens only when X and Y have the same sign
      but the result has the opposite sign.
    - We test the sign (MSB) of the 32-bit operands:
        acc_r[31]   : sign of accumulator (1 = negative, 0 = non-negative)
        prod32[31]  : sign of product extended to 32 bits
        sum[31]     : sign of result
      Positive overflow detected when both operands non-negative but result negative:
        pos_oflow = (~acc_r[31]) & (~prod32[31]) & (sum[31])
      Negative overflow detected when both operands negative but result non-negative:
        neg_oflow = (acc_r[31]) & (prod32[31]) & (~sum[31])

  Concrete numeric examples (illustrative)
    - Positive overflow:
        acc_r = 1_200_000_000  (sign=0)
        prod32 = 1_200_000_000 (sign=0)
        sum (32-bit two's complement) becomes negative -> pos_oflow = 1
    - Negative overflow:
        acc_r = -1_200_000_000 (sign=1)
        prod32 = -1_200_000_000 (sign=1)
        sum becomes positive -> neg_oflow = 1

  Safety / design note
    - Worst-case single product magnitude: 127 * 127 = 16129
    - For Tk = 64, worst-case sum magnitude = 64 * 16129 = 1,032,256 << 2^31
    - 32-bit accumulator is therefore sufficient for intended tiling; SAT still useful
      as defensive behaviour if tiles or accumulation depth change.

  Verification & DoD checklist
    - Unit tests (tb/unit/tb_mac8.sv) should include:
        * random vectors with multiple seeds (5 seeds required by DoD)
        * edge vectors that trigger pos/neg overflow
        * python golden dot-product checks for bit-exact behavior
    - Waveform (VCD/FSDB) snapshot saved for at least one overflow case.
*/

`ifndef MAC8_V
`define MAC8_V
`default_nettype none
// -----------------------------------------------------------------------------
// Title      : mac8
// File       : mac8.v
// Author     : Accel v1 Auto-Gen Assistant
// Description: Signed 8x8 -> 32-bit accumulate MAC with optional saturation.
//              Verilog-2001 compliant (no SystemVerilog keywords).
//
// Requirements Trace (examples):
//   REQ-ACCEL-MAC-01: Multiply two signed 8-bit operands each enabled cycle.
//   REQ-ACCEL-MAC-02: Accumulate product into signed 32-bit accumulator.
//   REQ-ACCEL-MAC-03: Provide synchronous clear (clr) and asynchronous reset.
//   REQ-ACCEL-MAC-04: Detect signed overflow and optionally saturate.
//   REQ-ACCEL-MAC-05: Provide sat_flag pulse when overflow occurs.
//   REQ-ACCEL-MAC-06: Deterministic hold when en=0.
//
// Safety / Notes:
//   Max product magnitude 127*127=16129; for K<=64 worst-case sum 1,032,256 < 2^31.
//   Saturation logic is defensive for future deeper accumulations.
// -----------------------------------------------------------------------------
// Parameters:
//   SAT (0/1) : 1 enables clamp to INT32_MIN/MAX on overflow; 0 allows wrap.
// -----------------------------------------------------------------------------
// Interface:
//   clk    : clock
//   rst_n  : async active-low reset
//   a,b    : signed 8-bit operands
//   clr    : sync clear (priority over en)
//   en     : accumulate enable
//   acc    : signed 32-bit accumulator output
//   sat_flag: 1-cycle pulse on overflow detection (even if SAT=0)
// -----------------------------------------------------------------------------
module mac8 #(parameter SAT = 0)(
    input  wire              clk,
    input  wire              rst_n,
    input  wire signed [7:0] a,
    input  wire signed [7:0] b,
    input  wire              clr,
    input  wire              en,
    output reg  signed [31:0] acc,
    output reg               sat_flag
);

    // Internal accumulator register
    reg signed [31:0] acc_r;
    reg               sat_r;
    wire signed [15:0] prod16 = a * b;      // 8x8 -> 16
    wire signed [31:0] prod32 = prod16;     // sign-extend to 32
    wire signed [31:0] sum = acc_r + prod32;
    wire pos_oflow = (~acc_r[31]) & (~prod32[31]) & (sum[31]);
    wire neg_oflow = (acc_r[31]) & (prod32[31]) & (~sum[31]);

    // Sequential logic
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            acc_r <= 32'sd0;  // Clear on reset
        end else if (clr) begin
            acc_r <= 32'sd0;  // Clear on command
        end else if (en) begin
            if (SAT && pos_oflow)
                acc_r <= 32'sh7FFFFFFF;
            else if (SAT && neg_oflow)
                acc_r <= 32'sh80000000;
            else
                acc_r <= sum;
        end else begin
            // hold
            acc_r <= acc_r;
            sat_r <= 1'b0;
        end
    end

    // Outputs
    always @(*) begin
        acc      = acc_r;
        sat_flag = sat_r;
    end

endmodule
`default_nettype wire
`endif
